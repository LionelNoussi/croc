module dma (
    ports
);
    
endmodule